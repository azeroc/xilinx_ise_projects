`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:19:45 01/16/2017 
// Design Name: 
// Module Name:    d_ff 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: Simple D-Flip-Flop
// 
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module d_ff(
    clk,
    d,
    q
);

input wire clk;
input wire d;
output reg q;

// Initialization
initial begin
    q = 0;
end

always@(posedge clk) begin
    q = d;
end

endmodule
